* SPICE 3f5 Level 8, Star-HSPICE Level 49, UTMOST Level 8

.lib cmos_models

* DATE: Feb 23/01

* LOT: T0BM WAF: 07

* Temperature_parameters=Default

.MODEL nmos NMOS ( LEVEL = 49

+VERSION = 3.1 TNOM = 27 TOX = 5.8E-9

+XJ = 1E-7 NCH = 2.3549E17 VTH0 = 0.3907535

+K1 = 0.4376003 K2 = 8.265151E-3 K3 = 4.214601E-3

+K3B = -3.7220937 W0 = 2.517345E-6 NLX = 2.310668E-7

+DVT0W = 0 DVT1W = 0 DVT2W = 0

+DVT0 = 0.2411602 DVT1 = 0.3707226 DVT2 = -0.5

+U0 = 316.5922683 UA = -9.89493E-10 UB = 2.154013E-18

+UC = 2.474632E-11 VSAT = 1.254499E5 A0 = 1.2735648

+AGS = 0.2428704 B0 = 2.579719E-8 B1 = -1E-7

+KETA = 4.87168E-4 A1 = 0 A2 = 0.5196633

+RDSW = 120 PRWG = 0.5 PRWB = -0.2

+WR = 1 WINT = 2.357855E-8 LINT = 1.210018E-9

+DWG = 2.292632E-9

+DWB = -9.94921E-10 VOFF = -0.1039771 NFACTOR = 1.3905578

+CIT = 0 CDSC = 2.4E-4 CDSCD = 0

+CDSCB = 0 ETA0 = 3.894977E-3 ETAB = 7.800632E-4

+DSUB = 0.0307944 PCLM = 1.7312397 PDIBLC1 = 0.999135

+PDIBLC2 = 4.850036E-3 PDIBLCB = -0.0866866 DROUT = 0.8612131

+PSCBE1 = 7.995844E10 PSCBE2 = 1.457011E-8 PVAG = 0.0099984

+DELTA = 0.01 RSH = 5 MOBMOD = 1

+PRT = 0 UTE = -1.5 KT1 = -0.11

+KT1L = 0 KT2 = 0.022 UA1 = 4.31E-9

+UB1 = -7.61E-18 UC1 = -5.6E-11 AT = 3.3E4

+WL = 0 WLN = 1 WW = -1.22182E-16

+WWN = 1.2127 WWL = 0 LL = 0

+LLN = 1 LW = 0 LWN = 1

+LWL = 0 CAPMOD = 2 XPART = 0.4

+CGDO = 3.11E-10 CGSO = 3.11E-10 CGBO = 1E-12

+CJ = 1.741905E-3 PB = 0.9876681 MJ = 0.4679558

+CJSW = 3.653429E-10 PBSW = 0.99 MJSW = 0.2943558

+CF = 0 PVTH0 = -0.01 PRDSW = 0

+PK2 = 2.589681E-3 WKETA = -1.866069E-3 LKETA = -0.0166961 )

*

.MODEL pmos PMOS ( LEVEL = 49

+VERSION = 3.1 TNOM = 27 TOX = 5.8E-9

+XJ = 1E-7 NCH = 4.1589E17 VTH0 = -0.583228

+K1 = 0.5999865 K2 = 6.150203E-3 K3 = 0

+K3B = 3.6314079 W0 = 1E-6 NLX = 1E-9

+DVT0W = 0 DVT1W = 0 DVT2W = 0

+DVT0 = 2.8749516 DVT1 = 0.7488605 DVT2 = -0.0917408

+U0 = 136.076212 UA = 2.023988E-9 UB = 1E-21

+UC = -9.26638E-11 VSAT = 2E5 A0 = 0.951197

+AGS = 0.20963 B0 = 1.345599E-6 B1 = 5E-6

+KETA = 0.0114727 A1 = 3.851541E-4 A2 = 0.614676

+RDSW = 1.496983E3 PRWG = -0.0440632 PRWB = -0.2945454

+WR = 1 WINT = 7.879211E-9 LINT = 2.894523E-8

+DWG = -1.112097E-8

+DWB = 9.815716E-9 VOFF = -0.1204623 NFACTOR = 1.2259401

+CIT = 0 CDSC = 2.4E-4 CDSCD = 0

+CDSCB = 0 ETA0 = 0.3325261 ETAB = -0.0623452

+DSUB = 0.9206875 PCLM = 0.833903 PDIBLC1 = 9.948506E-4

+PDIBLC2 = 0.0191187 PDIBLCB = -1E-3 DROUT = 0.9938581

+PSCBE1 = 2.887413E10 PSCBE2 = 8.325891E-9 PVAG = 0.8478443

+DELTA = 0.01 RSH = 3.6 MOBMOD = 1

+PRT = 0 UTE = -1.5 KT1 = -0.11

+KT1L = 0 KT2 = 0.022 UA1 = 4.31E-9

+UB1 = -7.61E-18 UC1 = -5.6E-11 AT = 3.3E4

+WL = 0 WLN = 1 WW = 0

+WWN = 1 WWL = 0 LL = 0

+LLN = 1 LW = 0 LWN = 1

+LWL = 0 CAPMOD = 2 XPART = 0.4

+CGDO = 2.68E-10 CGSO = 2.68E-10 CGBO = 1E-12

+CJ = 1.864957E-3 PB = 0.976468 MJ = 0.4614408

+CJSW = 3.118281E-10 PBSW = 0.6870843 MJSW = 0.3021929

+CF = 0 PVTH0 = 6.397941E-3 PRDSW = 30.410214

+PK2 = 2.100359E-3 WKETA = 5.428923E-3 LKETA = -0.0111599 )

*

.endl


